module rowRegularLight (CLOCK, RESET, PRELIGHT, LIGHTON);

	input CLOCK, RESET, PRELIGHT;
	output LIGHTON;
	
endmodule;