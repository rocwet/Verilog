/* NAME					|	thirtyTwoBitXor.sv
	-------------------------------------------------------------------------------------------------
	DESCRIPTION       |  determines if a is less than b
 ---------------------------------------------------------------------------------------------------
	PARAMETERS			|	TYPE					|	DESCRIPTION					
 ---------------------------------------------------------------------------------------------------
	outXOR		      |	OUTPUT [31:0]		|	Binary value if a is less than b (1 = true; 0 = false)
	A						|	INPUT  [31:0]		| 	input a
	B						|	INPUT  [31:0]		| 	input b
	#################################################################################################
	AUTHOR            | Minhhue H Khuu && Vivi Chuang
	ASSIGNMENT			| Lab 2: Register File
	CLASS					| EE 471
	DATE					| 02/17/2015
	#################################################################################################
*/ 
module thirtyTwoBitXor #(parameter WIDTH = 32)(outXOR, a, b); 
	output [WIDTH-1:0] outXOR; 
	input [WIDTH-1:0] a, b; 

	genvar i; 

	generate 
		for (i = 0; i < WIDTH; i++) begin: eachXOR
			xor x1 (outXOR[i], a[i], b[i]); //do we need "." infront ??
		end 
	endgenerate

endmodule


// testbench
module thirtyTwoBitXor_testbench();
	reg [31:0] a, b;

	wire [31:0] outXOR;

	thirtyTwoBitXor dut (.outXOR, .a, .b);

	 initial begin
		 #10 a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000000;
		 #10 a = 32'b00011111111110000000000000000000; b = 32'b00000000100000000000000000000000;
		 #10 a = 32'b00000000000000000000000000000001; b = 32'b10000000000000000000000000000000;
		 #10 a = 32'b00000000000000000000000000011000; b = 32'b00000000000000000000000000000001;
		 #10 a = 32'b10000000000000000000000000000000; b = 32'b00000000000000000111111111111111;
		 #10 a = 32'b10000000000000000000000000000001; b = 32'b00000000000000000001111111000000;
		 #10 a = 32'b00000000000000000000000000000000; b = 32'b11111111111111111111111111111111;
		 #10 a = 32'b00000000000000000001000000000000; b = 32'b00000000000000000000000000000000;
		 #10 a = 32'b00000000000000000000000000000000; b = 32'b00000000000000000000000000000100;

	 end 

endmodule 