module ccount(CLOCK, RESET, SW, OUT);
	input CLOCK, RESET;
	input [8:0] SW;
	output reg OUT;
	
	wire [19:0] ss;
	


		

endmodule